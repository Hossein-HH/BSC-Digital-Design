//* bitwise operations :
// ~(NOT), &(AND), |(OR), ^(XOR), ~^(XNOR)

//* logical :
// &&,||,!

//* shift : >>,<<

//* concatenation :
// {,}

//* assign
// نوشتن اساین برای مواقعی هست که بین یک خروجی و ورودی یک معادله
// همیشگی و ثابت وجود دارد
// assign A = ~B ;

//* always @(x or y or w)
// هر سيگنالي كه داخل اين بلاك قرار ميگيره و سمت چپ باشه
// بايد به عنوان متغير براي برنامه تعريف بشه
// reg با كمك

// سيگنال هاي ورودي يا اينپوت هيچ وقت نميتونن 
// reg 
// باشن

// در يك برنامه ميتونيم چندين
// always 
// بنويسيم كه هر كودوم با سيگنال هاي ورودي متفاوتي كار بكنن و اجرا بشن

//* case
// case(x)
// 0: command;
// 1: command;
// 2: command;
// endcase