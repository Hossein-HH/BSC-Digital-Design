module name
  // نوشتن اسم ماژول
  (
    // نوشتن خروجی ها
    doorOpen,
    //نوشتن ورودی ها
    doorSen
  );

  // خروجی

  output doorOpen;
  // نوشتن اسم خروجی ها

  reg doorOpen;
  // نوشتن اسم خروجی ها

  // متغیر چند بیتی
  // اگه نیاز به تعریف متغیر چند بیتی بود به این صورت مینویسیم
  // reg [3:0] a;
  // خط بالا تعریف یک متغیر 4 بیتی هست که با ارزش ترین بیت سمت چپ
  // قرار دارد

  // آرایه
  // اگه نیاز به تعریف آرایه بود به این صورت مینویسیم
  // reg a [3:0];
  // خط بالا تعریف یک آرایه 4 عنصری هست که هر عنصر 1 بیت دارد
  // وقتی میگوئیم 1 بیت دارد یعنی فقط 0 یا 1 میتوانیم
  // در آن قرار دهیم

  // آرایه ای از متغیر های چند بیتی
  // reg [3:0] a [5:0];
  // خط بالا تعریف یک آرایه با 6 عنصر هست که هر عنصر 4 بیت دارد

  // ورودی

  input doorSen;
  // نوشتن اسم ورودی ها



  always @(*)
    // در بلاک
    // always
    // شروطی که برای به وجود آمدن سیگنال های خروجی در صورت مسئله
    // داده میشود را اینجا مینویسیم

  begin
    // به عنوان مثال در خطوط زیر بررسی میشود که اگر مقدار سنسور درب
    // برابر با عدد 1 شده است درب را باز کند

    if (doorSen == 1)
    begin
      doorOpen = 1;
    end


  end
endmodule

////////////////////////////////

// تست بنچ

module name_tb;
  // نوشتن اسم ماژول تست بنچ و اضافه کردن
  // _tb
  //  به آخر اسم آن

  integer i;
  // تعریف متغیر برای حلقه ای که تست بنچ را تولید میکند از نوع اینتیجر

  // تعریف خروجی ها از نوع سیم یا همان
  // wire
  wire doorOpen;

  // تعریف خروجی ها از نوع متغیر یا همان
  // reg
  reg doorSen;

  // در اینجا نیز باید قبل از کلمه
  // uut
  // اسمی که برای ماژول اصلی انتخاب کردیم را بنوسیم
  // کوچک ترین اشتباه تایپی در این  قسمت منجر به عدم رسیدن به جواب میشود
  name uut(

         // نوشتن تابع
         // uut
         // جهت اتصال ماژول اصلی به تست بنچ

         // مقدار دهی نظیر به نظیر خروجی ها
         .doorOpen(doorOpen),
         // مقدار دهی نظیر به نظیر ورودی ها
         .doorSen(doorSen)
       );

  initial
    // نوشتن بلاک
    // initial
    // برای مقدار دادن به اینپوت ها یا همان ورودی های مسئله

  begin
    for (i = 0; i < 20; ++i)
      // یک حلقه به طول دلخواه (نه خیلی کم نه خیلی زیاد
      // (همین 20 یا 10 خوبه
    begin
      // برای تولید و ریختن آن در یک متغیر مشابه خط زیر عمل میکنیم
      // x = {$random} % 2;
      // برای تولید یک عدد تصادفی بین 
      // a,b => a < x < b
      // به صورت زیر عمل میکنیم
      // x = a + {$random} % b;
      // برای خط بالا فقط کافیست آ و بی را تغییر دهید
    end
  end
endmodule
